* Filtre RC passe-bas du premier ordre

* Parametres (alignes avec la DataFrame: R_val, C_val)
.param R_val = 1k
.param C_val = 100n

* Source d'entree : DC = 0, AC = 1 V
Vin in 0 0 AC 1

* Filtre RC : R en serie, C a la masse
R1 in out {R_val}
C1 out 0 {C_val}

* Balayage AC log : 1 Hz -> 1 MHz
.ac dec 100 1 1Meg

* Mesure de la frequence de coupure (-3 dB)
.meas ac fcut WHEN vdb(out) = -3

.end
