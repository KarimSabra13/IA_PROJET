* RC low-pass filter, first order

.param Rval = 1k
.param Cval = 100n

* Input source, AC amplitude 1 V
Vin in 0 AC 1

* R in series, C to ground
R1 in out {Rval}
C1 out 0 {Cval}

* AC sweep from 10 Hz to 1 MHz
.ac dec 100 10 1Meg

.end

